module module2()

reg [41:0] tab[0:39];
// reg[0:31] = value ; reg[32:36] = index of that value in table 1 ;reg[37:41] = index of that value in table 2; 

tab[0][0:31] =14; 
tab[0][32:36]=4;
tab[0][37:41]=18;
tab[1][0:31] =89; 
tab[1][32:36]=9;
tab[1][37:41]=9;
tab[2][0:31] =48; 
tab[2][32:36]=12;
tab[2][37:41]=8;
tab[3][0:31] =76; 
tab[3][32:36]=16;
tab[3][37:41]=16;
tab[4][0:31] =13; 
tab[4][32:36]=17;
tab[4][37:41]=5;
tab[5][0:31] =82; 
tab[5][32:36]=8;
tab[5][37:41]=2;
tab[6][0:31] =70; 
tab[6][32:36]=0;
tab[6][37:41]=10;
tab[7][0:31] =11; 
tab[7][32:36]=11;
tab[7][37:41]=19;
tab[8][0:31] =91; 
tab[8][32:36]=11;
tab[8][37:41]=11;
tab[9][0:31] =13; 
tab[9][32:36]=5;
tab[9][37:41]=17;
tab[10][0:31] =97; 
tab[10][32:36]=17;
tab[10][37:41]=13;


    
    
endmodule