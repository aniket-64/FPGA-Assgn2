module mod1 (
    output reg [31:0] table1 [19:0],
    output reg [31:0] table2 [19:0]
);

    table1[
    
endmodule