module module2();

    reg [31:0] val[0:39];
    reg [4:0] i1 [0:39];
    reg [4:0] i2 [0:39];
    reg cp [0:39];

val[0] =14; 
i1 [0]=4;
i2[0]=18;
cp[0]=1;
val[1] =89; 
i1[1]=9;
i2[1]=9;
    cp[1]=1;
val[2] =48; 
i1[2]=12;
i2[2]=8;
    cp[2]=1;
val[3] =76; 
i1[3]=16;
i2[3]=16;
    cp[3]=1;
val[4] =13; 
i1[4]=17;
i2[4]=5;
    cp[4]=1;
val[5]=82; 
i1[5]=8;
i2[5]=2;
    cp[5]=1;
val[6]=70; 
i1[6]=0;
i2[6]=10;
    cp[6]=1;
val[7]=11; 
i1[7]=11;
i2[7]=19;
    cp[7]=1;
val[8]=91; 
i1[8]=11;
i2[8]=11;
    cp[8]=1;
val[9] =13; 
i1[9]=5;
i2[9]=17;
    cp[9]=1;
val[10]=97; 
i1[10]=17;
i2[10]=13;
    cp[10]=1;


    
    
endmodule
